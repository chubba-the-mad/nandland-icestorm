module not_gate (
	input i_Switch_1,
	output o_LED_1);

assign o_LED_1 = ~i_Switch_1;

endmodule
